//`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08.05.2024 09:43:20
// Design Name: 
// Module Name: tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_maj_pca_score;
//Parameters
    parameter FP_SIZE = 64, PC_NUM = 5, MAJ_PC_NUM = 2;
    
// Inputs and Outputs

//********************************************************* USING 64 BIT BINARY *********************************************************************
//---------------------------------------------- CLOCK INSERTED ----------------------------------------------------------
 //   logic wire clk, reset,
//    reg [FP_SIZE-1:0] maj_eigen_values [0:MAJ_PC_NUM-1],
//    reg [FP_SIZE-1:0] maj_principal_comps [0:MAJ_PC_NUM-1],
//    reg [FP_SIZE-1:0] maj_pc_score
//------------------------------------------------------------------------------------------------------------------------
//---------------------------------------------- NO CLOCK INSERTED -------------------------------------------------------
//    reg [FP_SIZE-1:0] maj_eigen_values [0:MAJ_PC_NUM-1],
//    reg [FP_SIZE-1:0] maj_principal_comps [0:MAJ_PC_NUM-1],
//    reg [FP_SIZE-1:0] maj_pc_score
//------------------------------------------------------------------------------------------------------------------------
//***************************************************************************************************************************************************

//********************************************************* USING FLOATING POINT *********************************************************************
//---------------------------------------------- CLOCK INSERTED ----------------------------------------------------------
    logic clk, reset;
//    real maj_eigen_values [0:MAJ_PC_NUM-1];
//    real maj_principal_comps [0:MAJ_PC_NUM-1];
//    real maj_pc_score;
//------------------------------------------------------------------------------------------------------------------------
//---------------------------------------------- NO CLOCK INSERTED -------------------------------------------------------
    real maj_eigen_values [0:MAJ_PC_NUM-1];
    real maj_principal_comps [0:MAJ_PC_NUM-1];
    real maj_pc_score;
//------------------------------------------------------------------------------------------------------------------------
//***************************************************************************************************************************************************  
    
// Instantiaing the DUT
maj_pca_score
dut (
//---------------------------------------------- CLOCK ASSIGNMENTS ----------------------------------------------------------
//    .clk(clk), .reset(reset),
//------------------------------------------------------------------------------------------------------------------------
    .maj_eigen_values(maj_eigen_values),
    .maj_principal_comps(maj_principal_comps),
    .maj_pc_score(maj_pc_score)
);

initial begin
//---------------------------------------------- CLOCK ASSERTIONS ----------------------------------------------------------
$display($time, " << Starting the Simulation >>");
    reset = 1'b1;
    clk = 1'b1;

    #50 reset = ~reset;
////------------------------------------------------------------------------------------------------------------------------

//********************************************************* USING 64 BIT BINARY *********************************************************************

//***************************************************************************************************************************************************

//********************************************************* USING FLOATING POINT *********************************************************************
maj_eigen_values[0] =4;
maj_eigen_values[1] =3;

maj_principal_comps[0] = 2;
maj_principal_comps[1] = 3;
//***************************************************************************************************************************************************

end

    always begin
        #50 clk = ~clk; // Toggle the clock every 5 time units
    end

endmodule
