
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`include "pp_loop_interface.svh"
`include "pp_loop_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.values2Strm_U.if_read & AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.values2Strm_U.if_empty_n;
    assign fifo_intf_1.wr_en = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.values2Strm_U.if_write & AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.values2Strm_U.if_full_n;
    assign fifo_intf_1.fifo_rd_block = ~(AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.values2Strm_0_blk_n);
    assign fifo_intf_1.fifo_wr_block = ~(AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.values2Strm_0_blk_n);
    assign fifo_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.values2Strm_1_U.if_read & AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.values2Strm_1_U.if_empty_n;
    assign fifo_intf_2.wr_en = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.values2Strm_1_U.if_write & AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.values2Strm_1_U.if_full_n;
    assign fifo_intf_2.fifo_rd_block = ~(AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.values2Strm_1_blk_n);
    assign fifo_intf_2.fifo_wr_block = ~(AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.values2Strm_1_blk_n);
    assign fifo_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.rows_c_U.if_read & AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.rows_c_U.if_empty_n;
    assign fifo_intf_3.wr_en = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.rows_c_U.if_write & AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.rows_c_U.if_full_n;
    assign fifo_intf_3.fifo_rd_block = ~(AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.rows_blk_n);
    assign fifo_intf_3.fifo_wr_block = ~(AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.rows_c_blk_n);
    assign fifo_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.cols_c_U.if_read & AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.cols_c_U.if_empty_n;
    assign fifo_intf_4.wr_en = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.cols_c_U.if_write & AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.cols_c_U.if_full_n;
    assign fifo_intf_4.fifo_rd_block = ~(AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.cols_blk_n);
    assign fifo_intf_4.fifo_wr_block = ~(AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.cols_c_blk_n);
    assign fifo_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;

logic region_0_idle;
logic [31:0] region_0_start_cnt;
logic [31:0] region_0_done_cnt;
assign region_0_idle = (region_0_start_cnt == region_0_done_cnt) && AESL_inst_dut.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_start_cnt <= 32'h0;
    else if (AESL_inst_dut.ap_start == 1'b1 && AESL_inst_dut.ap_ready == 1'b1)
        region_0_start_cnt <= region_0_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_done_cnt <= 32'h0;
    else if (AESL_inst_dut.ap_done == 1'b1)
        region_0_done_cnt <= region_0_done_cnt + 32'h1;
    else;
end

logic region_1_idle;
logic [31:0] region_1_start_cnt;
logic [31:0] region_1_done_cnt;
assign region_1_idle = (region_1_start_cnt == region_1_done_cnt) && AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_1_start_cnt <= 32'h0;
    else if (AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.ap_start == 1'b1 && AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.ap_ready == 1'b1)
        region_1_start_cnt <= region_1_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_1_done_cnt <= 32'h0;
    else if (AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.ap_done == 1'b1 && AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.ap_continue == 1'b1)
        region_1_done_cnt <= region_1_done_cnt + 32'h1;
    else;
end


    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.real_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0 | ~AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.values2Strm_0_blk_n | ~AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.values2Strm_1_blk_n | ~AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.rows_c_blk_n | ~AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.cols_c_blk_n;
    assign process_intf_1.cin_stall = 1'b0;
    assign process_intf_1.cout_stall = 1'b0;
    assign process_intf_1.region_idle = region_1_idle;
    assign process_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_start;
    assign process_intf_2.pin_stall = 1'b0 | ~AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.rows_blk_n | ~AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.cols_blk_n | ~AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.values2Strm_0_blk_n | ~AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.values2Strm_1_blk_n;
    assign process_intf_2.pout_stall = 1'b0;
    assign process_intf_2.cin_stall = 1'b0;
    assign process_intf_2.cout_stall = 1'b0;
    assign process_intf_2.region_idle = region_1_idle;
    assign process_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_dut.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_dut.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_dut.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.ap_done;
    assign module_intf_6.ap_continue = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.ap_continue;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_dut.grp_implement_fu_147.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_dut.grp_implement_fu_147.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_dut.grp_implement_fu_147.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = 1'b0;
    assign module_intf_19.ap_ready = 1'b0;
    assign module_intf_19.ap_done = 1'b0;
    assign module_intf_19.ap_continue = 1'b0;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_start;
    assign module_intf_30.ap_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_ready;
    assign module_intf_30.ap_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_done;
    assign module_intf_30.ap_continue = 1'b1;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_start;
    assign module_intf_31.ap_ready = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_ready;
    assign module_intf_31.ap_done = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_done;
    assign module_intf_31.ap_continue = 1'b1;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;

    pp_loop_intf #(4) pp_loop_intf_1(clock,reset);
    assign pp_loop_intf_1.pre_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_ST_fsm_state1;
    assign pp_loop_intf_1.pre_states_valid = 1'b1;
    assign pp_loop_intf_1.post_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_ST_fsm_state9;
    assign pp_loop_intf_1.post_states_valid[0] = 1'b1;
    assign pp_loop_intf_1.post_loop_state1 = 4'h0;
    assign pp_loop_intf_1.post_states_valid[1] = 1'b0;
    assign pp_loop_intf_1.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_1.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_enable_reg_pp0_iter6;
    assign pp_loop_intf_1.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.loop_quit_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.quit_at_end = 1'b1;
    assign pp_loop_intf_1.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.ap_CS_fsm;
    assign pp_loop_intf_1.finish = finish;
    csv_file_dump pp_loop_csv_dumper_1;
    pp_loop_monitor #(4) pp_loop_monitor_1;
    pp_loop_intf #(6) pp_loop_intf_2(clock,reset);
    assign pp_loop_intf_2.pre_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_ST_fsm_state1;
    assign pp_loop_intf_2.pre_states_valid = 1'b1;
    assign pp_loop_intf_2.post_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_ST_fsm_state5;
    assign pp_loop_intf_2.post_states_valid[0] = 1'b1;
    assign pp_loop_intf_2.post_loop_state1 = 6'h0;
    assign pp_loop_intf_2.post_states_valid[1] = 1'b0;
    assign pp_loop_intf_2.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_2.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_2.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_2.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_2.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_2.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_2.loop_quit_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_2.quit_at_end = 1'b1;
    assign pp_loop_intf_2.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.ap_CS_fsm;
    assign pp_loop_intf_2.finish = finish;
    csv_file_dump pp_loop_csv_dumper_2;
    pp_loop_monitor #(6) pp_loop_monitor_2;
    pp_loop_intf #(7) pp_loop_intf_3(clock,reset);
    assign pp_loop_intf_3.pre_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_ST_fsm_state1;
    assign pp_loop_intf_3.pre_states_valid = 1'b1;
    assign pp_loop_intf_3.post_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_ST_fsm_state7;
    assign pp_loop_intf_3.post_states_valid[0] = 1'b1;
    assign pp_loop_intf_3.post_loop_state1 = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_ST_fsm_state8;
    assign pp_loop_intf_3.post_states_valid[1] = 1'b1;
    assign pp_loop_intf_3.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_3.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_3.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_3.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_3.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_enable_reg_pp0_iter1;
    assign pp_loop_intf_3.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_3.loop_quit_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_ST_fsm_pp0_stage3;
    assign pp_loop_intf_3.quit_at_end = 1'b0;
    assign pp_loop_intf_3.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_125_1_fu_297.ap_CS_fsm;
    assign pp_loop_intf_3.finish = finish;
    csv_file_dump pp_loop_csv_dumper_3;
    pp_loop_monitor #(7) pp_loop_monitor_3;
    seq_loop_intf#(82) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.ap_ST_fsm_state36;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.ap_ST_fsm_state1;
    assign seq_loop_intf_1.post_states_valid = 1'b1;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.ap_ST_fsm_state37;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.ap_ST_fsm_state37;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.ap_ST_fsm_state82;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(82) seq_loop_monitor_1;
    seq_loop_intf#(5) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_2.post_states_valid = 1'b1;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(5) seq_loop_monitor_2;
    seq_loop_intf#(5) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_3.pre_states_valid = 1'b1;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_3.post_states_valid = 1'b1;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(5) seq_loop_monitor_3;
    seq_loop_intf#(39) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_ST_fsm_state37;
    assign seq_loop_intf_4.pre_states_valid = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_4.post_states_valid = 1'b1;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_ST_fsm_state38;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_ST_fsm_state38;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.ap_ST_fsm_state39;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(39) seq_loop_monitor_4;
    seq_loop_intf#(21) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_dut.grp_implement_fu_147.ap_ST_fsm_state6;
    assign seq_loop_intf_5.pre_states_valid = 1'b1;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_dut.grp_implement_fu_147.ap_ST_fsm_state13;
    assign seq_loop_intf_5.post_states_valid = 1'b1;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_dut.grp_implement_fu_147.ap_ST_fsm_state7;
    assign seq_loop_intf_5.quit_states_valid = 1'b1;
    assign seq_loop_intf_5.cur_state = AESL_inst_dut.grp_implement_fu_147.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_dut.grp_implement_fu_147.ap_ST_fsm_state7;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_dut.grp_implement_fu_147.ap_ST_fsm_state12;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(21) seq_loop_monitor_5;
    seq_loop_intf#(21) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state3;
    assign seq_loop_intf_6.pre_states_valid = 1'b1;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state14;
    assign seq_loop_intf_6.post_states_valid = 1'b1;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state4;
    assign seq_loop_intf_6.quit_states_valid = 1'b1;
    assign seq_loop_intf_6.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state4;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state13;
    assign seq_loop_intf_6.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(21) seq_loop_monitor_6;
    seq_loop_intf#(21) seq_loop_intf_7(clock,reset);
    assign seq_loop_intf_7.pre_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state14;
    assign seq_loop_intf_7.pre_states_valid = 1'b1;
    assign seq_loop_intf_7.post_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state14;
    assign seq_loop_intf_7.post_states_valid = 1'b1;
    assign seq_loop_intf_7.quit_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state15;
    assign seq_loop_intf_7.quit_states_valid = 1'b1;
    assign seq_loop_intf_7.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_CS_fsm;
    assign seq_loop_intf_7.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state15;
    assign seq_loop_intf_7.iter_end_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state21;
    assign seq_loop_intf_7.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_7.one_state_loop = 1'b0;
    assign seq_loop_intf_7.one_state_block = 1'b0;
    assign seq_loop_intf_7.finish = finish;
    csv_file_dump seq_loop_csv_dumper_7;
    seq_loop_monitor #(21) seq_loop_monitor_7;
    seq_loop_intf#(21) seq_loop_intf_8(clock,reset);
    assign seq_loop_intf_8.pre_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state4;
    assign seq_loop_intf_8.pre_states_valid = 1'b1;
    assign seq_loop_intf_8.post_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state1;
    assign seq_loop_intf_8.post_states_valid = 1'b1;
    assign seq_loop_intf_8.quit_loop_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state14;
    assign seq_loop_intf_8.quit_states_valid = 1'b1;
    assign seq_loop_intf_8.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_CS_fsm;
    assign seq_loop_intf_8.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state14;
    assign seq_loop_intf_8.iter_end_state0 = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.ap_ST_fsm_state15;
    assign seq_loop_intf_8.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_8.one_state_loop = 1'b0;
    assign seq_loop_intf_8.one_state_block = 1'b0;
    assign seq_loop_intf_8.finish = finish;
    csv_file_dump seq_loop_csv_dumper_8;
    seq_loop_monitor #(21) seq_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_ST_fsm_state1;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_ST_fsm_state1;
    assign upc_loop_intf_1.quit_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_ST_fsm_state1;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_1.quit_block = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_1.iter_start_enable = 1'b1;
    assign upc_loop_intf_1.iter_end_enable = 1'b1;
    assign upc_loop_intf_1.quit_enable = 1'b1;
    assign upc_loop_intf_1.loop_start = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_VITIS_LOOP_283_1_fu_368.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_2.quit_enable = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_2.loop_start = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a1_fu_376.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;
    upc_loop_intf#(2) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_3.quit_state = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_enable_reg_pp0_iter5;
    assign upc_loop_intf_3.quit_enable = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_enable_reg_pp0_iter5;
    assign upc_loop_intf_3.loop_start = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_dut.grp_aveImpl_double_15_80_1_2_16_s_fu_119.grp_aveImpl_double_15_80_1_2_16_Pipeline_loop_a2_fu_389.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(2) upc_loop_monitor_3;
    upc_loop_intf#(2) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_4.quit_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_enable_reg_pp0_iter9;
    assign upc_loop_intf_4.quit_enable = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_enable_reg_pp0_iter9;
    assign upc_loop_intf_4.loop_start = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart1_double_15_80_1_2_16_U0.grp_covCorePart1_double_15_80_1_2_16_Pipeline_loop_c2_fu_153.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(2) upc_loop_monitor_4;
    upc_loop_intf#(16) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_ST_fsm_pp0_stage4;
    assign upc_loop_intf_5.quit_state = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_ST_fsm_pp0_stage4;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_block_pp0_stage4_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_block_pp0_stage4_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_enable_reg_pp0_iter9;
    assign upc_loop_intf_5.quit_enable = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_enable_reg_pp0_iter9;
    assign upc_loop_intf_5.loop_start = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_dut.grp_covCoreWrapper_double_15_80_1_2_16_s_fu_129.covCorePart2_double_15_2_16_U0.grp_covCorePart2_double_15_2_16_Pipeline_VITIS_LOOP_245_2_fu_80.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(16) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_6.quit_enable = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_6.loop_start = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_277_1_VITIS_LOOP_278_2_fu_138.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b1;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_7.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_7.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_init_A_VITIS_LOOP_91_1_fu_267.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b1;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_ST_fsm_state1;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_ST_fsm_state1;
    assign upc_loop_intf_8.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_ST_fsm_state1;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_8.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_8.iter_start_enable = 1'b1;
    assign upc_loop_intf_8.iter_end_enable = 1'b1;
    assign upc_loop_intf_8.quit_enable = 1'b1;
    assign upc_loop_intf_8.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_142_1_fu_313.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b1;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_9.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_9.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_precal_fu_320.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_cal_fu_328.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(1) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_enable_reg_pp0_iter6;
    assign upc_loop_intf_11.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_enable_reg_pp0_iter6;
    assign upc_loop_intf_11.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_VITIS_LOOP_1005_1_fu_336.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(1) upc_loop_monitor_11;
    upc_loop_intf#(2) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_enable_reg_pp0_iter69;
    assign upc_loop_intf_12.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_enable_reg_pp0_iter69;
    assign upc_loop_intf_12.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_Jacobi_svd_double_16_1_16_Pipeline_Loop_jacobi2x2_fu_348.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b1;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(2) upc_loop_monitor_12;
    upc_loop_intf#(4) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_13.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_enable_reg_pp0_iter6;
    assign upc_loop_intf_13.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_enable_reg_pp0_iter6;
    assign upc_loop_intf_13.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollRow_double_16_1_16_9_fu_401.ap_done_int;
    assign upc_loop_intf_13.loop_continue = 1'b1;
    assign upc_loop_intf_13.quit_at_end = 1'b1;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(4) upc_loop_monitor_13;
    upc_loop_intf#(4) upc_loop_intf_14(clock,reset);
    assign upc_loop_intf_14.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_CS_fsm;
    assign upc_loop_intf_14.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_14.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_14.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_14.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_14.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_14.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_enable_reg_pp0_iter6;
    assign upc_loop_intf_14.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_enable_reg_pp0_iter6;
    assign upc_loop_intf_14.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_start;
    assign upc_loop_intf_14.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_ready;
    assign upc_loop_intf_14.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_gesvdj_2D_double_16_1_16_s_fu_280.grp_Jacobi_svd_double_16_1_16_s_fu_85.grp_funcDataflow_double_16_1_16_8_fu_390.grp_unrollCol_double_16_1_16_10_fu_412.ap_done_int;
    assign upc_loop_intf_14.loop_continue = 1'b1;
    assign upc_loop_intf_14.quit_at_end = 1'b1;
    assign upc_loop_intf_14.finish = finish;
    csv_file_dump upc_loop_csv_dumper_14;
    upc_loop_monitor #(4) upc_loop_monitor_14;
    upc_loop_intf#(1) upc_loop_intf_15(clock,reset);
    assign upc_loop_intf_15.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_CS_fsm;
    assign upc_loop_intf_15.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_15.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_15.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_15.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_start;
    assign upc_loop_intf_15.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_ready;
    assign upc_loop_intf_15.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_Loop_postcal_VITIS_LOOP_113_2_fu_287.ap_done_int;
    assign upc_loop_intf_15.loop_continue = 1'b1;
    assign upc_loop_intf_15.quit_at_end = 1'b1;
    assign upc_loop_intf_15.finish = finish;
    csv_file_dump upc_loop_csv_dumper_15;
    upc_loop_monitor #(1) upc_loop_monitor_15;
    upc_loop_intf#(1) upc_loop_intf_16(clock,reset);
    assign upc_loop_intf_16.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_CS_fsm;
    assign upc_loop_intf_16.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_16.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_16.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_start;
    assign upc_loop_intf_16.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_ready;
    assign upc_loop_intf_16.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop_fu_308.ap_done_int;
    assign upc_loop_intf_16.loop_continue = 1'b1;
    assign upc_loop_intf_16.quit_at_end = 1'b1;
    assign upc_loop_intf_16.finish = finish;
    csv_file_dump upc_loop_csv_dumper_16;
    upc_loop_monitor #(1) upc_loop_monitor_16;
    upc_loop_intf#(1) upc_loop_intf_17(clock,reset);
    assign upc_loop_intf_17.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_CS_fsm;
    assign upc_loop_intf_17.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_17.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_17.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_start;
    assign upc_loop_intf_17.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_ready;
    assign upc_loop_intf_17.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_NSort_shift_buf_Loop12_fu_314.ap_done_int;
    assign upc_loop_intf_17.loop_continue = 1'b1;
    assign upc_loop_intf_17.quit_at_end = 1'b1;
    assign upc_loop_intf_17.finish = finish;
    csv_file_dump upc_loop_csv_dumper_17;
    upc_loop_monitor #(1) upc_loop_monitor_17;
    upc_loop_intf#(1) upc_loop_intf_18(clock,reset);
    assign upc_loop_intf_18.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_CS_fsm;
    assign upc_loop_intf_18.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_18.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_enable_reg_pp0_iter37;
    assign upc_loop_intf_18.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_enable_reg_pp0_iter37;
    assign upc_loop_intf_18.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_start;
    assign upc_loop_intf_18.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_ready;
    assign upc_loop_intf_18.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_filtermat_loop_VITIS_LOOP_160_1_fu_320.ap_done_int;
    assign upc_loop_intf_18.loop_continue = 1'b1;
    assign upc_loop_intf_18.quit_at_end = 1'b1;
    assign upc_loop_intf_18.finish = finish;
    csv_file_dump upc_loop_csv_dumper_18;
    upc_loop_monitor #(1) upc_loop_monitor_18;
    upc_loop_intf#(1) upc_loop_intf_19(clock,reset);
    assign upc_loop_intf_19.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_CS_fsm;
    assign upc_loop_intf_19.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_19.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_enable_reg_pp0_iter38;
    assign upc_loop_intf_19.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_enable_reg_pp0_iter38;
    assign upc_loop_intf_19.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_start;
    assign upc_loop_intf_19.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_ready;
    assign upc_loop_intf_19.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_PCA_Sign_Normalization_Loop_VITIS_LOOP_214_1_fu_335.ap_done_int;
    assign upc_loop_intf_19.loop_continue = 1'b1;
    assign upc_loop_intf_19.quit_at_end = 1'b1;
    assign upc_loop_intf_19.finish = finish;
    csv_file_dump upc_loop_csv_dumper_19;
    upc_loop_monitor #(1) upc_loop_monitor_19;
    upc_loop_intf#(1) upc_loop_intf_20(clock,reset);
    assign upc_loop_intf_20.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_CS_fsm;
    assign upc_loop_intf_20.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_ST_fsm_state1;
    assign upc_loop_intf_20.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_ST_fsm_state1;
    assign upc_loop_intf_20.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_ST_fsm_state1;
    assign upc_loop_intf_20.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_20.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_20.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_20.iter_start_enable = 1'b1;
    assign upc_loop_intf_20.iter_end_enable = 1'b1;
    assign upc_loop_intf_20.quit_enable = 1'b1;
    assign upc_loop_intf_20.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_start;
    assign upc_loop_intf_20.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_ready;
    assign upc_loop_intf_20.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_238_2_fu_349.ap_done_int;
    assign upc_loop_intf_20.loop_continue = 1'b1;
    assign upc_loop_intf_20.quit_at_end = 1'b1;
    assign upc_loop_intf_20.finish = finish;
    csv_file_dump upc_loop_csv_dumper_20;
    upc_loop_monitor #(1) upc_loop_monitor_20;
    upc_loop_intf#(1) upc_loop_intf_21(clock,reset);
    assign upc_loop_intf_21.cur_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_CS_fsm;
    assign upc_loop_intf_21.iter_start_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_end_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.quit_state = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_start_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_end_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.quit_block = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_start_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_21.iter_end_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_21.quit_enable = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_21.loop_start = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_start;
    assign upc_loop_intf_21.loop_ready = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_ready;
    assign upc_loop_intf_21.loop_done = AESL_inst_dut.grp_implement_fu_147.grp_implement_Pipeline_VITIS_LOOP_244_4_fu_360.ap_done_int;
    assign upc_loop_intf_21.loop_continue = 1'b1;
    assign upc_loop_intf_21.quit_at_end = 1'b1;
    assign upc_loop_intf_21.finish = finish;
    csv_file_dump upc_loop_csv_dumper_21;
    upc_loop_monitor #(1) upc_loop_monitor_21;
    upc_loop_intf#(1) upc_loop_intf_22(clock,reset);
    assign upc_loop_intf_22.cur_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_CS_fsm;
    assign upc_loop_intf_22.iter_start_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_end_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.quit_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_start_block = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_end_block = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.quit_block = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_start_enable = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_22.iter_end_enable = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_enable_reg_pp0_iter12;
    assign upc_loop_intf_22.quit_enable = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_enable_reg_pp0_iter12;
    assign upc_loop_intf_22.loop_start = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_start;
    assign upc_loop_intf_22.loop_ready = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_ready;
    assign upc_loop_intf_22.loop_done = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_350_2_VITIS_LOOP_351_3_fu_156.ap_done_int;
    assign upc_loop_intf_22.loop_continue = 1'b1;
    assign upc_loop_intf_22.quit_at_end = 1'b1;
    assign upc_loop_intf_22.finish = finish;
    csv_file_dump upc_loop_csv_dumper_22;
    upc_loop_monitor #(1) upc_loop_monitor_22;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);

    pp_loop_csv_dumper_1 = new("./pp_loop_status1.csv");
    pp_loop_monitor_1 = new(pp_loop_intf_1,pp_loop_csv_dumper_1);
    pp_loop_csv_dumper_2 = new("./pp_loop_status2.csv");
    pp_loop_monitor_2 = new(pp_loop_intf_2,pp_loop_csv_dumper_2);
    pp_loop_csv_dumper_3 = new("./pp_loop_status3.csv");
    pp_loop_monitor_3 = new(pp_loop_intf_3,pp_loop_csv_dumper_3);


    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);
    seq_loop_csv_dumper_7 = new("./seq_loop_status7.csv");
    seq_loop_monitor_7 = new(seq_loop_intf_7,seq_loop_csv_dumper_7);
    seq_loop_csv_dumper_8 = new("./seq_loop_status8.csv");
    seq_loop_monitor_8 = new(seq_loop_intf_8,seq_loop_csv_dumper_8);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);
    upc_loop_csv_dumper_14 = new("./upc_loop_status14.csv");
    upc_loop_monitor_14 = new(upc_loop_intf_14,upc_loop_csv_dumper_14);
    upc_loop_csv_dumper_15 = new("./upc_loop_status15.csv");
    upc_loop_monitor_15 = new(upc_loop_intf_15,upc_loop_csv_dumper_15);
    upc_loop_csv_dumper_16 = new("./upc_loop_status16.csv");
    upc_loop_monitor_16 = new(upc_loop_intf_16,upc_loop_csv_dumper_16);
    upc_loop_csv_dumper_17 = new("./upc_loop_status17.csv");
    upc_loop_monitor_17 = new(upc_loop_intf_17,upc_loop_csv_dumper_17);
    upc_loop_csv_dumper_18 = new("./upc_loop_status18.csv");
    upc_loop_monitor_18 = new(upc_loop_intf_18,upc_loop_csv_dumper_18);
    upc_loop_csv_dumper_19 = new("./upc_loop_status19.csv");
    upc_loop_monitor_19 = new(upc_loop_intf_19,upc_loop_csv_dumper_19);
    upc_loop_csv_dumper_20 = new("./upc_loop_status20.csv");
    upc_loop_monitor_20 = new(upc_loop_intf_20,upc_loop_csv_dumper_20);
    upc_loop_csv_dumper_21 = new("./upc_loop_status21.csv");
    upc_loop_monitor_21 = new(upc_loop_intf_21,upc_loop_csv_dumper_21);
    upc_loop_csv_dumper_22 = new("./upc_loop_status22.csv");
    upc_loop_monitor_22 = new(upc_loop_intf_22,upc_loop_csv_dumper_22);

    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_1);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_2);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_7);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_15);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_16);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_17);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_18);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_19);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_20);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_21);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_22);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1 || deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
