////`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////////
//// Company: 
//// Engineer: 
//// 
//// Create Date: 08.05.2024 09:43:20
//// Design Name: 
//// Module Name: tb
//// Project Name: 
//// Target Devices: 
//// Tool Versions: 
//// Description: 
//// 
//// Dependencies: 
//// 
//// Revision:
//// Revision 0.01 - File Created
//// Additional Comments:
//// 
////////////////////////////////////////////////////////////////////////////////////


//module tb_maj_dot;
////Parameters
//    parameter FP_SIZE = 64, PC_NUM = 5, MAJ_PC_NUM = 2;
    
//// Inputs and Outputs
////********************************************************* USING 64 BIT BINARY *********************************************************************
////---------------------------------------------- CLOCK INSERTED ----------------------------------------------------------
// //   logic clk, reset;
////    reg [FP_SIZE-1:0] common_vector [0:PC_NUM -1];
////    reg [FP_SIZE-1:0] long_vector [0:MAJ_PC_NUM-1][0:PC_NUM -1];
////    logic [FP_SIZE-1:0] out_vector [0:MAJ_PC_NUM-1];
////------------------------------------------------------------------------------------------------------------------------
////---------------------------------------------- NO CLOCK INSERTED -------------------------------------------------------
////    reg [FP_SIZE-1:0] common_vector [0:PC_NUM -1];
////    reg [FP_SIZE-1:0] long_vector [0:MAJ_PC_NUM-1][0:PC_NUM -1];
////    logic [FP_SIZE-1:0] out_vector [0:MAJ_PC_NUM-1];
////------------------------------------------------------------------------------------------------------------------------

////***************************************************************************************************************************************************

////********************************************************* USING FLOATING POINT *********************************************************************

////---------------------------------------------- CLOCK INSERTED ----------------------------------------------------------
//    logic clk, reset;
////    real common_vector [0:PC_NUM -1];
////    real long_vector [0:MAJ_PC_NUM-1][0:PC_NUM -1];
////    real out_vector [0:MAJ_PC_NUM-1];
////------------------------------------------------------------------------------------------------------------------------
////---------------------------------------------- NO CLOCK INSERTED -------------------------------------------------------
//    real common_vector [0:PC_NUM -1];
//    real long_vector [0:MAJ_PC_NUM-1][0:PC_NUM -1];
//    real out_vector [0:MAJ_PC_NUM-1];
////------------------------------------------------------------------------------------------------------------------------
////***************************************************************************************************************************************************  
    
//// Instantiaing the DUT
//maj_dot
//dut (
////---------------------------------------------- CLOCK ASSIGNMENTS ----------------------------------------------------------
////    .clk(clk), .reset(reset),
////------------------------------------------------------------------------------------------------------------------------
//    .common_vector(common_vector),
//    .long_vector(long_vector),
//    .out_vector(out_vector)
//);



//initial begin

////---------------------------------------------- CLOCK ASSERTIONS ----------------------------------------------------------
//$display($time, " << Starting the Simulation >>");
//    reset = 1'b1;
//    clk = 1'b1;

//    #50 reset = ~reset;
//////------------------------------------------------------------------------------------------------------------------------

////********************************************************* USING 64 BIT BINARY *********************************************************************
////common_vector[0] = 64'b0100000000001000000000000000000000000000000000000000000000000000;
////common_vector[1] = 64'b0100000000010000000000000000000000000000000000000000000000000000;
////common_vector[2] = 64'b0100000000000000000000000000000000000000000000000000000000000000;
////common_vector[3] = 64'b0100000000010100000000000000000000000000000000000000000000000000;
////common_vector[4] = 64'b0011111111110000000000000000000000000000000000000000000000000000;


////long_vector[0][0] = 64'b0100000000001000000000000000000000000000000000000000000000000000;
////long_vector[0][1] = 64'b0100000000000000000000000000000000000000000000000000000000000000;
////long_vector[0][2] = 64'b0011111111110000000000000000000000000000000000000000000000000000;
////long_vector[0][3] = 64'b0100000000100000000000000000000000000000000000000000000000000000;
////long_vector[0][4] = 64'b0100000000010100000000000000000000000000000000000000000000000000;

////long_vector[1][0] = 64'b0011111111110000000000000000000000000000000000000000000000000000;
////long_vector[1][1] = 64'b0011111111110000000000000000000000000000000000000000000000000000;
////long_vector[1][2] = 64'b0011111111110000000000000000000000000000000000000000000000000000;
////long_vector[1][3] = 64'b0011111111110000000000000000000000000000000000000000000000000000;
////long_vector[1][4] = 64'b0011111111110000000000000000000000000000000000000000000000000000;
////***************************************************************************************************************************************************

////********************************************************* USING FLOATING POINT *********************************************************************
//common_vector[0] = 3;
//common_vector[1] = 4;
//common_vector[2] = 2;
//common_vector[3] = 5;
//common_vector[4] = 1;


//long_vector[0][0] = 3;
//long_vector[0][1] = 2;
//long_vector[0][2] = 1;
//long_vector[0][3] = 8;
//long_vector[0][4] = 5;

//long_vector[1][0] = 1;
//long_vector[1][1] = 1;
//long_vector[1][2] = 1;
//long_vector[1][3] = 1;
//long_vector[1][4] = 1;
////***************************************************************************************************************************************************


////#100; // Specify a runtime of 100 ps
//end

//    always begin
//        #50 clk = ~clk; // Toggle the clock every 5 time units
//    end


//endmodule
