//`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08.05.2024 09:43:20
// Design Name: 
// Module Name: tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_threshold_compare;
//Parameters
    parameter FP_SIZE = 64, PC_NUM = 5, MAJ_PC_NUM = 2;
    
// Inputs and Outputs
//********************************************************* USING 64 BIT BINARY *********************************************************************
//---------------------------------------------- CLOCK INSERTED ----------------------------------------------------------
 //   logic clk, reset;
//    reg [FP_SIZE-1:0] common_vector [0:PC_NUM -1];
//    reg [FP_SIZE-1:0] long_vector [0:MAJ_PC_NUM-1][0:PC_NUM -1];
//    logic [FP_SIZE-1:0] out_vector [0:MAJ_PC_NUM-1];
//------------------------------------------------------------------------------------------------------------------------
//---------------------------------------------- NO CLOCK INSERTED -------------------------------------------------------
//    reg [FP_SIZE-1:0] common_vector [0:PC_NUM -1];
//    reg [FP_SIZE-1:0] long_vector [0:MAJ_PC_NUM-1][0:PC_NUM -1];
//    logic [FP_SIZE-1:0] out_vector [0:MAJ_PC_NUM-1];
//------------------------------------------------------------------------------------------------------------------------

//***************************************************************************************************************************************************

//********************************************************* USING FLOATING POINT *********************************************************************

//---------------------------------------------- CLOCK INSERTED ----------------------------------------------------------
    logic clk, reset;
//    real common_vector [0:PC_NUM -1];
//    real long_vector [0:MAJ_PC_NUM-1][0:PC_NUM -1];
//    real out_vector [0:MAJ_PC_NUM-1];
//------------------------------------------------------------------------------------------------------------------------
//---------------------------------------------- NO CLOCK INSERTED -------------------------------------------------------
    real maj_pc_score;
    real min_pc_score;
    real out_d;

//------------------------------------------------------------------------------------------------------------------------
//***************************************************************************************************************************************************  
    
// Instantiaing the DUT
threshold_compare
dut (
//---------------------------------------------- CLOCK ASSIGNMENTS ----------------------------------------------------------
//    .clk(clk), .reset(reset),
//------------------------------------------------------------------------------------------------------------------------
    .maj_pc_score(maj_pc_score),
    .min_pc_score(min_pc_score),
    .out_d(out_d)
);



initial begin

//---------------------------------------------- CLOCK ASSERTIONS ----------------------------------------------------------
$display($time, " << Starting the Simulation >>");
    reset = 1'b1;
    clk = 1'b1;

    #50 reset = ~reset;
////------------------------------------------------------------------------------------------------------------------------

//********************************************************* USING 64 BIT BINARY *********************************************************************

//***************************************************************************************************************************************************

//********************************************************* USING FLOATING POINT *********************************************************************
//t_max = 7.364668875,
//t_min = 18.48677496

//~~~~~~~~~~~~ Both Higher~~~~~~~~~~~
//    maj_pc_score = 8.13231;
//    min_pc_score = 20.34534;
    
   
////~~~~~~~~~~~~ Only Maj Higher ~~~~~~~~~~~
//    maj_pc_score = 11.1231234;
//    min_pc_score = 5.2452456;
    
//    //~~~~~~~~~~~~ Only Min Higher ~~~~~~~~~~~
//    maj_pc_score = 4.2545151;
//    min_pc_score = 32.545341;
    
//    //~~~~~~~~~~~~ Both Lower~~~~~~~~~~~
    maj_pc_score = 3.2341134;
    min_pc_score = 6.2546566;
//***************************************************************************************************************************************************


//#100; // Specify a runtime of 100 ps
end

    always begin
        #50 clk = ~clk; // Toggle the clock every 5 time units
    end


endmodule
